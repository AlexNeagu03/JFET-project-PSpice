* D:\Desktop\TEMA DE CASA DE\wroklab1\Schematic2TEMA.sch

* Schematics Version 9.1 - Web Update 1
* Tue Jan 17 14:38:13 2023



** Analysis setup **
.DC LIN V_VCC 0 25 1 
+ LIN V_VGS 0 3 1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2TEMA.net"
.INC "Schematic2TEMA.als"


.probe


.END
